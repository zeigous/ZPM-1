
module FetchBuffer(
    input clk,
    input clkEn,
    input rst
);
    
endmodule
