
module FetchEngine(
    input clk,
    input clkEn,
    input rst

);

    
endmodule : FetchEngine