
module L1ICache(
    input clk,
    input clkEn,
    input rst
);

endmodule
