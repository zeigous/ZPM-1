module core(
    input clk,
    input clkEn,
    input rst
);
    
endmodule : core
